library verilog;
use verilog.vl_types.all;
entity pratica2 is
    port(
        clock           : in     vl_logic;
        ir              : in     vl_logic_vector(8 downto 0);
        din             : in     vl_logic_vector(15 downto 0);
        run             : in     vl_logic;
        resetn          : in     vl_logic;
        q               : out    vl_logic_vector(15 downto 0);
        r0t             : out    vl_logic_vector(15 downto 0);
        r1t             : out    vl_logic_vector(15 downto 0);
        r2t             : out    vl_logic_vector(15 downto 0);
        r3t             : out    vl_logic_vector(15 downto 0);
        r4t             : out    vl_logic_vector(15 downto 0);
        r5t             : out    vl_logic_vector(15 downto 0);
        r6t             : out    vl_logic_vector(15 downto 0);
        r7t             : out    vl_logic_vector(15 downto 0);
        At              : out    vl_logic_vector(15 downto 0);
        Gt              : out    vl_logic_vector(15 downto 0);
        r0_int          : out    vl_logic;
        r1_int          : out    vl_logic;
        r2_int          : out    vl_logic;
        r3_int          : out    vl_logic;
        r4_int          : out    vl_logic;
        r5_int          : out    vl_logic;
        r6_int          : out    vl_logic;
        r7_int          : out    vl_logic;
        r0_outt         : out    vl_logic;
        r1_outt         : out    vl_logic;
        r2_outt         : out    vl_logic;
        r3_outt         : out    vl_logic;
        r4_outt         : out    vl_logic;
        r5_outt         : out    vl_logic;
        r6_outt         : out    vl_logic;
        r7_outt         : out    vl_logic;
        g_outt          : out    vl_logic;
        dinoutt         : out    vl_logic;
        a_int           : out    vl_logic;
        g_int           : out    vl_logic;
        add_subt        : out    vl_logic;
        donet           : out    vl_logic;
        addsub_outt     : out    vl_logic_vector(15 downto 0);
        buswiret        : out    vl_logic_vector(15 downto 0)
    );
end pratica2;
